
B0 7 10 23 jjSFQ1 area=40
B1 8 12 24 jjSFQ1 area=40
B2 7 14 25 jjSFQ1 area=40
B3 8 16 26 jjSFQ1 area=40
B4 20 21 27 jjSFQ1 area=40
B5 20 22 28 jjSFQ1 area=40
I0 0 6 pwl(0 0 0.1ns 0 0.19ns 10u)
I1 0 7 pwl(0 0 0.09n 0 0.1n Ide )
I2 0 8 pwl(0 0 0.09n 0 0.1n 73u)
I3 0 20 pwl(0 0 0.09n 0 0.1n 73u)
K1 L11 L10 1
K2 L15 L14 1
K3 L6 L7 1
K4 L4 L5 1
L0 6 9 100n
L1 7 11 50n
L2 8 2 57.5p
L3 6 13 100n
L4 9 4 250p
L5 10 0 20p
L6 11 15 200p
L7 12 0 20p
L8 2 17 0p
L9 14 0 20p
L10 16 0 20p
L11 19 18 20p
L12 20 19 57.5p
L13 21 0 20p
L14 22 0 20p
L15 0 5 20p
R0 1 0 1
R1 0 3 1
R2 13 0 R=v(3)+1e-6
R3 15 0 R=v(1)+0.0502
R4 17 5 R=v(1)+1.55e-3
R5 0 4 R=v(1)+4.008
R6 18 0 R=v(1)+1.55e-3
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)
V1 3 0 pwl(0 0 4.999n 0 5n 5e3 5.2n 5e3 5.201n 0)

.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
