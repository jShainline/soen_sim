
B0 5 6 13 jjSFQ1 area=40
B1 5 7 14 jjSFQ1 area=40
B2 10 11 15 jjSFQ1 area=40
B3 10 12 16 jjSFQ1 area=40
I0 0 4 pwl(0 0 1ns 0 101ns 17u)
I1 0 5 pwl(0 0 0.09n 0 0.1n Ide )
I2 0 10 pwl(0 0 0.09n 0 0.1n 73u)
K1 L4 L3 1
K2 L8 L7 1
K3 L1 L2 1
L0 5 2 57.5p
L1 4 0 200p
L2 6 0 20p
L3 7 0 20p
L4 9 8 20p
L5 10 9 57.5p
L6 11 0 20p
L7 12 0 20p
L8 0 3 20p
R0 1 0 1
R1 2 3 R=v(1)+1.55e-3
R2 8 0 R=v(1)+1.55e-3
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)

.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
