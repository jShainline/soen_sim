
B0 5 13 25 jjSFQ1 area=40
B1 10 17 26 jjSFQ1 area=40
B2 5 19 27 jjSFQ1 area=40
B3 6 0 28 jjSFQ1 area=40
B4 7 0 29 jjSFQ1 area=40
B5 10 23 30 jjSFQ1 area=40
B6 11 0 31 jjSFQ1 area=40
B7 12 0 32 jjSFQ1 area=40
B8 21 0 33 jjSFQ2 area=40
I0 0 5 pwl(0 0 0.09n 0 0.1n 76u)
I1 0 6 pwl(0 0 0.09n 0 0.1ns 36u)
I2 0 7 pwl(0 0 0.09n 0 0.1ns 35u)
I3 0 8 pwl(0 0 0.09n 0 0.1n 35u)
I4 0 9 pwl(0 0 0.1ns 0 0.19ns 10u)
I5 0 10 pwl(0 0 0.09n 0 0.1n 72u)
I6 0 11 pwl(0 0 0.09n 0 0.1ns 36u)
I7 0 12 pwl(0 0 0.09n 0 0.1ns 35u)
K1 L17 L15 1
K2 L9 L10 -1
K3 L14 L8 1
K4 L12 L13 1
L0 5 6 200p
L1 6 7 77.5p
L2 7 14 7.75n
L3 8 15 1f
L4 9 16 100n
L5 10 11 200p
L6 11 12 77.5p
L7 12 18 50n
L8 13 0 20p
L9 14 20 200p
L10 8 21 20p
L11 9 22 100n
L12 16 4 250p
L13 17 0 20p
L14 18 24 200p
L15 19 0 20p
L16 23 0 20p
L17 2 0 20p
R0 1 0 1
R1 15 2 R=v(1)+1e-3
R2 0 3 1
R3 24 0 R=v(1)+0.1004
R4 20 0 R=v(1)+0.0195
R5 22 0 R=v(3)+1e-6
R6 0 4 R=v(1)+4.005
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)
V1 3 0 pwl(0 0 4.999n 0 5n 5e3 5.2n 5e3 5.201n 0)
.model jjSFQ2 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 0f, vshunt=0.25mV)

*hysteretic JJ for driving xTron
.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
.save @I5[c]
.save @I2[c]
.save @I4[c]
.save @I6[c]
.save @I7[c]
.save @I0[c]
.save @I1[c]
.save @I3[c]
