
B0 4 7 11 jjSFQ1 area=40
B1 4 8 12 jjSFQ1 area=40
B2 5 9 13 jjSFQ1 area=40
B3 6 10 14 jjSFQ1 area=40
I0 0 3 pwl(0 0 1ns 0 101ns 18u)
 I1 0 4 pwl(0 0 0.09n 0 0.1n 81u )
I2 0 5 pwl(0 0 0.09n 0 0.1ns 15u)
I3 0 6 pwl(0 0 0.09n 0 0.1ns 25u)
K1 L3 L4 1
L0 4 5 65p
L1 5 6 65p
L2 6 2 65p
L3 3 0 200p
L4 7 0 20p
L5 8 0 20p
L6 9 0 1f
L7 10 0 1f
R0 1 0 1
R1 2 0 R=v(1)+1.3e-3
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)

.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
.control
set maxdata=2560000
tran 1p 101n
write ./ne_4jj_direct_drive_lin_ramp_alt_ind_Ldrv200pH_Lnr20pH20pH_Ide81.00uA_taunf50.00ns_dt01.0ps.dat L2#branch L3#branch
quit
.endc
