
B0 2 6 11 jjSFQ1 area=40
B1 2 7 12 jjSFQ1 area=40
B2 2 8 13 jjSFQ1 area=40
 I0 0 2 pwl(0 0 0.2ns 0 0.3ns  85.00u )
 I1 0 9 pwl(0 0 0.4ns 0 0.5ns  2.471534u )
 I2 0 10 pwl(0 0 0.6ns 0 0.7ns 10.669522u )
K1 L2 L3 1
K2 L4 L5 1
L0 3 2 77.5n
L1 3 4 200p
L2 9 0 200p
 L3 6 0 35.00p 
L4 10 0 400p
L5 7 5 12.5p
L6 8 5 12.5p
L7 5 0 1f
R0 1 0 1
R1 4 0 R=v(1)+1e-6
V0 1 0 pwl(0 1e6 0.9ns 1e6 1ns 0)
.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
.control
set maxdata=2560000
tran 1p 20.300000n
write ./dend_3jj_nest_cnst_drv_seek_rt_arry_Ib085.00uA_Lp35.00pH_Ip02.471534uA_Iex10.669522.dat i(L1) v(2) v(13)
quit
.endc
