
B0 4 11 22 jjSFQ1 area=40
B1 8 14 23 jjSFQ1 area=40
B2 4 16 24 jjSFQ1 area=40
B3 5 17 25 jjSFQ1 area=40
B4 6 18 26 jjSFQ1 area=40
B5 8 20 27 jjSFQ1 area=40
B6 9 0 28 jjSFQ1 area=40
B7 10 0 29 jjSFQ1 area=40
 I0 0 4 pwl(0 0 0.09n 0 0.1n 82u )
I1 0 5 pwl(0 0 0.09n 0 0.1ns 15u)
I2 0 6 pwl(0 0 0.09n 0 0.1ns 25u)
I3 0 7 pwl(0 0 0.1ns 0 0.19ns 10u)
 I4 0 8 pwl(0 0 0.09n 0 0.1n 78u )
I5 0 9 pwl(0 0 0.09n 0 0.1ns 36u)
I6 0 10 pwl(0 0 0.09n 0 0.1ns 35u)
K1 L11 L7 1
K2 L9 L10 1
L0 4 5 65p
L1 5 6 65p
L2 6 12 65p
L3 7 13 100n
L4 8 9 200p
L5 9 10 77.5p
L6 10 15 50n 
L7 11 0 20p
L8 7 19 100n
L9 13 3 250p
L10 14 0 20p
L11 15 21 200p
L12 16 0 20p
L13 17 0 1f
L14 18 0 1f
L15 20 0 20p
R0 1 0 1
R1 12 0 R=v(1)+1.56e-3
R2 0 2 1
 R3 21 0 R=v(1)+0.1 
R4 19 0 R=v(2)+1e-6
R5 0 3 R=v(1)+4.005
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)
V1 2 0 pwl(0 0 4.999n 0 5n 5e3 5.2n 5e3 5.201n 0)

.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
.control
set maxdata=2560000
tran 10p 300n
write ./ne_4jj_1pls_Isy78.00uA_Ide82.00uA_tausi0500.00ns.dat L9#branch L11#branch L2#branch
quit
.endc
