 
B0 3 4 7 jjSFQ1 area=40
B1 3 6 8 jjSFQ1 area=40
I0 0 2 pwl(0 0 0.09ns 0 0.1ns Idrive )
I1 0 3 pwl(0 0 0.09n 0 0.1n Ide )
K1 L1 L2 1
L0 3 5 77.5p
L1 2 0 200p
L2 4 0 20p
L3 6 0 20p
R0 1 0 1
R1 5 0 R=v(1)+1.55e-3
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)

.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
