
B0 4 7 9 jjSFQ1 area=40
B1 4 8 10 jjSFQ1 area=40
B2 5 0 11 jjSFQ1 area=40
B3 6 0 12 jjSFQ1 area=40
 I0 0 3 pwl(0 0 0.1ns 0 0.19ns 13.85u )
 I1 0 4 pwl(0 0 0.09n 0 0.1n 68.0u )
I2 0 5 pwl(0 0 0.09n 0 0.1ns 32u)
I3 0 6 pwl(0 0 0.09n 0 0.1ns 35u)
K1 L3 L4 1
L0 4 5 77.5p
L1 5 6 77.5p
L2 6 2 77.5p
L3 3 0 200p
L4 7 0 20p
L5 8 0 20p
R0 1 0 1
R1 2 0 R=v(1)+1.55e-3
V0 1 0 pwl(0 1e5 0.2ns 1e5 0.3ns 0)
.model jjSFQ1 jj(rtype=0, cct=1, vg=2.8m, icrit=1u, cap= 5f, vshunt=0.25mV)
.save @I2[c]
.save @I1[c]
.save @I3[c]
.save @I0[c]
.control
set maxdata=2560000
tran 1p 250n
write ./ne_4jj_direct_drive_cnst_drv_Lnr20pH20pH_Ide68.00uA_Ldrv200pH_Idrv13.85_taunf50.00ns_dt01.0ps.dat L2#branch
quit
.endc
